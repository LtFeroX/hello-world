include IEEE
